library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- TODO: Add libraries.

entity template is
  generic (
    -- TODO: Add generics.
  );
  port (
    -- TODO: Add ports.
  );
end;

architecture rtl of template is

  -- TODO: Add signals.

begin
  
  combinational : process () -- Add ports.
  begin
    -- TODO: Add combinational logic.
  end process;

  -- TODO: Add properties.
  -- Properties:
  -- skip psl default clock is rising_edge(clk);

end;

